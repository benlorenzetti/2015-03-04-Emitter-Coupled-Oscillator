*** simple.cir ***
* Nodes:
* cc, ee, c1, b1, e1, c2, b2, e2

Vcc cc gnd dc 24V ac 0V
Vee ee gnd dc 0V ac 0V
Rc1 cc c1 98.6
Rc2 cc c2 98.2
Q1 c1 b1 e1 model1
Q2 c2 b2 e2 model2
Re1 e1 ee 899
Re2 e2 ee 899
Rb1 b1 c2 147.8
Rb3 b2 c1 146.5
Rb2 b1 ee 1791
Rb4 b2 ee 1796
Cc e1 e2 50.4E-12


* .model <name> <type> (par1=value1 par2=value2 ...)
* VAF = forward Early voltage
* BF = forward beta; forward common-emitter gain
* CJE = base-emitter zero-bias junction capacitance
* CJC = base-collector zero-bias junction capacitance
* TS = transport saturation current
* NF = forward mode ideality factor

.model model1 npn (BF=176 CJC=3.291p CJE=5.255p IS=1E-16 VAF=121 NF=1)
.model model2 npn (BF=153 CJC=3.199p CJE=5.235p IS=1E-16 VAF=120 NF=1)

.control
set filetype=ascii
* tran <tstep> <tstop> <tstart> <tmax> ; the last two are optional

tran 1E-10 1E-6 1E-10
plot v(c1)
write simple-transient.txt v(c1)

tran 1E-10 101E-7 100E-7 1E-10
plot v(c1) v(c2) 
plot v(e1)-v(e2)


